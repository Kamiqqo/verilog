assign atan_table[00] = 32'b00100000000000000000000000000000; // atan(2^0)
assign atan_table[01] = 32'b00010010111001000000010100011101; // atan(2^-1)
assign atan_table[02] = 32'b00001001111110110011100001011011; // atan(2^-2)
assign atan_table[03] = 32'b00000101000100010001000111010100; // atan(2^-3) 
assign atan_table[04] = 32'b00000010100010110000110101000011; // atan(2^-4)
assign atan_table[05] = 32'b00000001010001011101011111100001; // atan(2^-5)
assign atan_table[06] = 32'b00000000101000101111011000011110; // atan(2^-6)
assign atan_table[07] = 32'b00000000010100010111110001010101; // atan(2^-7)
assign atan_table[08] = 32'b00000000001010001011111001010011; // atan(2^-8)
assign atan_table[09] = 32'b00000000000101000101111100101110; // atan(2^-9)
assign atan_table[10] = 32'b00000000000010100010111110011000; // atan(2^-10)
assign atan_table[11] = 32'b00000000000001010001011111001100; // atan(2^-11)
assign atan_table[12] = 32'b00000000000000101000101111100110; // atan(2^-12)
assign atan_table[13] = 32'b00000000000000010100010111110011; // atan(2^-13)
assign atan_table[14] = 32'b00000000000000001010001011111001; // atan(2^-14)
assign atan_table[15] = 32'b00000000000000000101000101111101; // atan(2^-15)
assign atan_table[16] = 32'b00000000000000000010100010111110; // atan(2^-16)
assign atan_table[17] = 32'b00000000000000000001010001011111; // atan(2^-17)
assign atan_table[18] = 32'b00000000000000000000101000101111; // atan(2^-18)
assign atan_table[19] = 32'b00000000000000000000010100011000; // atan(2^-19)
assign atan_table[20] = 32'b00000000000000000000001010001100; // atan(2^-20)
assign atan_table[21] = 32'b00000000000000000000000101000110; // atan(2^-21)
assign atan_table[22] = 32'b00000000000000000000000010100011; // atan(2^-22)
assign atan_table[23] = 32'b00000000000000000000000001010001; // atan(2^-23)
assign atan_table[24] = 32'b00000000000000000000000000101000; // atan(2^-24)
assign atan_table[25] = 32'b00000000000000000000000000010100; // atan(2^-25)
assign atan_table[26] = 32'b00000000000000000000000000001010; // atan(2^-26)
assign atan_table[27] = 32'b00000000000000000000000000000101; // atan(2^-27)
assign atan_table[28] = 32'b00000000000000000000000000000010; // atan(2^-28)
assign atan_table[29] = 32'b00000000000000000000000000000001; // atan(2^-29)
assign atan_table[30] = 32'b00000000000000000000000000000000; // atan(2^-30)
